VERSION 5.8 ;

MACRO greyhound_logo
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN tt_logo 0 0 ;
  SIZE 450.0 BY 450.0 ;

  OBS
    LAYER TopMetal2 ;
      RECT 0 0 450.0 450.0 ;
  END
END greyhound_logo
