`default_nettype none

module greyhound_logo ();
endmodule
